module PS2_keyboardController()
	
	
	
endmodule
