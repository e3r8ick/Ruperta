module ProcesadorARM()

endmodule
